# JSXE Swedish properties file
# $Id$
# Currently maintained by Patrik Johansson <patjoh@itstud.chalmers.se>
#:mode=properties:
#:tabSize=4:indentSize=4:noTabs=true:
#:folding=explicit:collapseFolds=1:

#{{{ common properties

common.ok=OK
common.cancel=Avbryt
common.close=StÃ¤ng
common.apply=VerkstÃ¤ll
common.more=Mer
common.insert=Infoga
common.add=LÃ¤gg till
common.remove=Ta bort
common.moveUp=Flytta upp
common.moveDown=Flytta ner
common.cut=Klipp ut
common.copy=Kopiera
common.paste=Klistra in
common.find=SÃ¶k...
common.findnext=SÃ¶k nÃ¤sta

#}}}

#{{{ Global Options
global.options.title=Globala instÃ¤llningar
#}}}

#{{{ File Menu Items
File.New=Ny
File.Open=Ã–ppna...
File.Recent=Senaste filer
File.Save=Spara
File.SaveAs=Spara som...
File.Reload=LÃ¤s om
File.Recent=Senaste filer
File.Close=StÃ¤ng
File.CloseAll=StÃ¤ng alla
File.Exit=Avsluta
#}}}

Tools.Options=InstÃ¤llningar...
Tools.Plugin=Hanterare fÃ¶r insticksprogram...
Plugin.Manager.Title=Hanterare fÃ¶r insticksprogram
Help.About=Om jsXe...
