# JSXE tree view Swedish properties file
# $Id$
# Currently maintained by Patrik Johansson <patjoh@itstud.chalmers.se>
#:mode=properties:
#:tabSize=4:indentSize=4:noTabs=true:
#:folding=explicit:collapseFolds=1:

TreeView.RenameNode=Ta bort nod
TreeView.RemoveNode=Ta bort nod
TreeView.AddAttribute=Lägg till attribut
TreeView.RemoveAttribute=Ta bort attribut
TreeView.EditNode=Redigera nod
