# JSXE Swedish properties file
# $Id$
# Currently maintained by Patrik Johansson <patjoh@itstud.chalmers.se>
#:mode=properties:
#:tabSize=4:indentSize=4:noTabs=true:
#:folding=explicit:collapseFolds=1:

SourceView.Cut=Klipp ut
SourceView.Copy=Kopiera
SourceView.Paste=Klistra in
SourceView.Find=Sök...
SourceView.FindNext=Sök nästa
