# JSXE Swedish properties file
# $Id$
# Currently maintained by Patrik Johansson <patjoh@itstud.chalmers.se>
#:mode=properties:
#:tabSize=4:indentSize=4:noTabs=true:
#:folding=explicit:collapseFolds=1:

#{{{ common properties

common.ok=OK
common.cancel=Avbryt
common.close=Stäng
common.apply=Verkställ
common.more=Mer
common.insert=Infoga
common.add=Lägg till
common.remove=Ta bort
common.moveUp=Flytta upp
common.moveDown=Flytta ner

#}}}

#{{{ Global Options
global.options.title=Globala inställningar
#}}}

#{{{ File Menu Items
File.New=Ny
File.Open=Öppna...
File.Recent=Senaste filer
File.Save=Spara
File.SaveAs=Spara som...
File.Reload=Läs om
File.Recent=Senaste filer
File.Close=Stäng
File.CloseAll=Stäng alla
File.Exit=Avsluta
#}}}

Edit.Node.Dialog.Title=Redigera nod
View.Tree=Trädvy
View.Source=Källkodsvy
Tools.Options=Inställningar...
Tools.Plugin=Hanterare för insticksprogram...
Plugin.Manager.Title=Hanterare för insticksprogram
Help.About=Om jsXe...

